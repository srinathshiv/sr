library ieee;
use ieee.std_logic_1164.all;

entity sr is
port (
    
);
end sr;

architecture rtrl of sr is


begin

end rtl;
